/***********************************************************************\
| Module:              bit_synchronizer
| Author:              Alex Hare
| Last Updated:        01/29/2021
| Function:            Synchronizes to when a packet is recieved. Will
|                      detect incoming packets
| Inputs:              
| Output:              
| Additional comments: Largely based on Benson, B. "Design of a Low-Cost 
|                      Underwater Acoustic Modem for Short-Range Sensor 
|                      Networks", UC San Diego, 2010
\***********************************************************************/
module set_threshold();

endmodule
